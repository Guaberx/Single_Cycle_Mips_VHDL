library ieee;
use ieee.std_logic_1164.all;

package muxes is
	
	type mux_32 is array (natural range <>) of std_logic_vector;

end package;