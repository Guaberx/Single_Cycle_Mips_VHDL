library verilog;
use verilog.vl_types.all;
entity monociclo_vlg_vec_tst is
end monociclo_vlg_vec_tst;
